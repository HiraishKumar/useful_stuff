module calc_diff(
    input signed [31:0] learn_in;
    input signed [127:0] grad_in;
    output signed [31:0] step_size
);



    
endmodule